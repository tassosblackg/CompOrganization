----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    18:54:35 03/17/2015 
-- Design Name: 
-- Module Name:    PC - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PC is
    Port ( addressIn : in  STD_LOGIC_vector(31 downto 0);
           LdEn : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           reset : in  STD_LOGIC;
           addressOut : out  STD_LOGIC_vector(31 downto 0));
end PC;

architecture Behavioral of PC is

begin
	process(clk)
	begin
	if clk'event and clk='1' then
	if reset='1' then
	addressOut<="00000000000000000000000000000000";
	elsif LdEn='1' then
	addressOut<=addressIn;
	end if;
	end if;
	end process;

end Behavioral;
